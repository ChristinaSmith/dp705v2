// Generator.bsv
// Copyright (c) 2012 Atomic Rules LLC - ALL RIGHTS RESERVED
// Christina Smith

import GetPut     ::*;
import FIFO       ::*;
import Vector     ::*;
import tbDefs     ::*;

interface Generatorv2Ifc;
  interface Get#(Mesg) src;
endinterface

module mkGeneratorv2(Generatorv2Ifc);

// state instanced here
FIFO#(Mesg)                  mesgOutF   <- mkFIFO;
Reg#(Bit#(8))                count      <- mkReg(0);
Reg#(Vector#(4, Bit#(8)))    patternV   <- mkReg(unpack('h00010203));
Reg#(Bit#(8))                mesgLen    <- mkReg(40);
Reg#(Vector#(4, Bit#(8)))    initV      <- mkReg(unpack('h01020304));
Reg#(Bool)                   tmp        <- mkReg(True);

function Bit#(8) addFour (Bit#(8) x) = x + 4;
function Bit#(8) addOne  (Bit#(8) x) = x + 1;

// rules here
rule genMesg;
  if(count < mesgLen) begin
    mesgOutF.enq(tagged ValidNotEOP pack(patternV));
    patternV <= map(addFour, patternV);
    count <= count + 1;
  end
  else if(count == mesgLen) begin
    mesgOutF.enq(tagged ValidEOP pack(patternV));
    patternV <= initV;
    initV <= map(addOne, initV);
    $display("genMesg2");
  end
endrule

//rule genEOP(count == mesgLen);
//  mesgOutF.enq(tagged ValidEOP pack(patternV));
//  patternV <= initV;
//  initV <= map(addOne, initV);
//endrule

//rule gobble;
//  $display("%0x",mesgOutF.first);
//  mesgOutF.deq;
//endrule

// interfaces provided here
interface src = toGet(mesgOutF);
endmodule
